module EvenPipe(clk, reset);
	input	clk, reset;
	
endmodule